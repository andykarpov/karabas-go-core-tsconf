/*
 * Copyright (c) 2013, Stefan Kristiansson <stefan.kristiansson@saunalahti.fi>
 * All rights reserved.
 *
 * Redistribution and use in source and non-source forms, with or without
 * modification, are permitted provided that the following conditions are met:
 *     * Redistributions of source code must retain the above copyright
 *       notice, this list of conditions and the following disclaimer.
 *     * Redistributions in non-source form must reproduce the above copyright
 *       notice, this list of conditions and the following disclaimer in the
 *       documentation and/or other materials provided with the distribution.
 *
 * THIS WORK IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
 * AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
 * THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR
 * PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
 * CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,
 * EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO,
 * PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
 * LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
 * ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
 * (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
 * WORK, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
 */

module i2s_rx #(
	parameter AUDIO_DW		= 16
)(
   input wire         clk,
	input	wire			sclk,
	input	wire			rst,

	input	wire			lrclk,
	input	wire			sdata,

	// Parallel datastreams
	output reg [AUDIO_DW-1:0]	left_chan,
	output reg [AUDIO_DW-1:0]	right_chan
);

reg [AUDIO_DW-1:0]	left;
reg [AUDIO_DW-1:0]	right;
reg			lrclk_r;
wire			lrclk_nedge;

assign lrclk_nedge = !lrclk & lrclk_r;

always @(posedge sclk)
	lrclk_r <= lrclk;

// sdata msb is valid one clock cycle after lrclk switches
always @(posedge sclk)
	if (lrclk_r)
		right <= {right[AUDIO_DW-2:0], sdata};
	else
		left <= {left[AUDIO_DW-2:0], sdata};

reg [AUDIO_DW-1:0] left_chan_r, right_chan_r;
reg rdy;
always @(posedge sclk) begin
	rdy <= 1'b0;
	if (rst) begin
		left_chan_r <= 0;
		right_chan_r <= 0;
	end else if (lrclk_nedge) begin
		rdy <= 1'b1;
		left_chan_r <= left;
		right_chan_r <= {right[AUDIO_DW-2:0], sdata};
	end
end

// transfer rdy
reg [1:0] rdy_r;
always @(posedge clk)
	rdy_r <= {rdy_r[0], rdy};

// transfer audio into clk domain
always @(posedge clk) begin
	if (rdy_r == 2'b10) begin // falling edge
	    left_chan <= left_chan_r;
	    right_chan <= right_chan_r;
	end
end


endmodule
