////////////////////////////////////////////////////////////////////////////////
//
//  PS2-to-Kempston Mouse v2
//  (C) 2017,2018 Sorgelig
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//
////////////////////////////////////////////////////////////////////////////////

module kempston_mouse
(
	input wire clk,
	input wire reset,

	input wire [7:0] ms_x,
	input wire [7:0] ms_y,
	input wire [3:0] ms_z,
	input wire [2:0] ms_b,
	input wire ms_upd,

	input wire [2:0] addr,
	output wire sel,
	output wire [7:0] dout
);

assign dout = data;
assign sel  = port_sel;

reg [11:0] dx;
reg [11:0] dy;
reg  [3:0] dz;

reg  [7:0] data;
reg        port_sel;

always @* begin
	port_sel = 1;
	casex(addr)
		 3'b011: data = dx[7:0];
		 3'b111: data = dy[7:0];
		 3'bX10: data = {dz, 1'b1, ~ms_b[2:0]};
		default: {port_sel,data} = 8'hFF;
	endcase
end

reg old_status;
always @(posedge clk) begin
	old_status <= ms_upd;

	if(reset) begin
		dx <= 128; // dx != dy for better mouse detection
		dy <= 0;
		dz <= 4'b1111;
	end
	else if(old_status != ms_upd) begin
		dx <= dx + ms_x;
		dy <= dy - ms_y;
		dz <= dz - ms_z;
	end
end

endmodule
