`timescale 1ns / 1ps
`default_nettype none

/*
 HDMI PLL chain to produce a pixelclock as well as x5 clock pair for hdmi serializer based on 
 detected frequency from the input clock clk.
 If the measured clk frequency is 28 MHz, then the clk_ref (28 MHz) will be passed directly to 5x PLL,
 otherwise the reconfigurable DCM_CLKGEN will be programmed and used via 8MHz base clock clk_8.
 The clk_8 clock will be multiplied to 3...10 to produce a desired 24...80MHz clock.
*/

module hdmi_pll(
	input wire clk, // muxed 28 from TS or 24...80 from FT (to measure only)
	input wire clk_ref, // 28 reference clock
	input wire clk_8, // 8 MHz clock (generated by design as base clock for FT812)
	input wire reset,
	input wire vdac2_sel, // selected ft source
	output wire clk_hdmi, // x5
	output wire clk_hdmi_n, // x5 180deg
	output wire clk_pix, // x1
	output wire clk_pix2, // x1/2
	output wire [7:0] freq, // detected frequency 28,24,32,40,56,64,72,80Mhz
	output wire locked,
	output wire o_reset
);

// freq counter
wire [7:0] hdmi_freq;
freq_counter freq_counter_inst(
	.i_clk_ref(clk_ref),
	.i_vdac2_sel(vdac2_sel),
	.i_clk_test(clk),
	.i_reset(reset),
	.o_freq(hdmi_freq)
);
assign freq = prev_hdmi_freq;

// detect freq change
reg hdmi_reset;
reg [7:0] prev_hdmi_freq;
reg prev_vdac2_sel;
always @(posedge clk_ref)
begin
	hdmi_reset <= 1'b0;
	// reset when switching back to 28 mhz
	if (~vdac2_sel && prev_vdac2_sel != vdac2_sel) begin
		hdmi_reset <= 1'b1;
	end
	// reset to reconfigure dcm
	else if (vdac2_sel && prog_done) begin
		if (prev_hdmi_freq != hdmi_freq) hdmi_reset <= 1'b1;
		prev_hdmi_freq <= hdmi_freq;
	end
	prev_vdac2_sel <= vdac2_sel;
end

// programming data for dcm_clkgen
reg [15:0] fctl; // {M,D}
reg [24:0] prog_data, prog_en;
always @(posedge clk_ref) begin
	if (hdmi_reset) begin
		case (hdmi_freq)
			8'd24: fctl <= {16'd3, 16'd1}; // M 3, D 1
			8'd32: fctl <= {16'd4, 16'd1}; // M 4, D 1
			8'd40: fctl <= {16'd5, 16'd1}; // M 5, D 1
			8'd48: fctl <= {16'd6, 16'd1}; // M 6, D 1
			8'd56: fctl <= {16'd7, 16'd1}; // M 7, D 1
			8'd64: fctl <= {16'd8, 16'd1}; // M 8, D 1
			8'd72: fctl <= {16'd9, 16'd1}; // M 9, D 1
			8'd80: fctl <= {16'd10, 16'd1}; // M 10, D 1		
			default: fctl <= {16'd10, 16'd1}; // M 10, D 1
		endcase
	end
end

// following https://docs.amd.com/v/u/en-US/ug382 section Dynamic Frequency Synthesis
always @(posedge clk_ref) begin
	if (hdmi_reset) begin
		// serial prog_data[0] : 10 - loadD command, D[0:7], 00 - gap, 11 - loadM command, M[0:7], 00 - gap, 1 - go.
		// serial prog_en[0]   : 11,               11111111, 00 - gap, 11,               11111111, 00 - gap, 0 - go.
		prog_data <= {1'b0, 2'b00, fctl[15:8]-1, 2'b11, 2'b00, fctl[7:0]-1, 2'b01};
		prog_en <=   {1'b1, 2'b00, 8'b11111111,  2'b11, 2'b00, 8'b11111111, 2'b11}; 
	end else begin
		prog_en   <= { 1'b0, prog_en  [24:1] };
		prog_data <= { 1'b0, prog_data[24:1] };
	end
end

// reconfigurable dcm to multiply and divide the clkin to a programmed M and D values
wire clkgen, prog_done, locked_dcm;
DCM_CLKGEN
  #(.CLKFXDV_DIVIDE        (2),
    .CLKFX_DIVIDE          (1),
    .CLKFX_MULTIPLY        (10), 
    .SPREAD_SPECTRUM       ("NONE"),
    .STARTUP_WAIT          ("FALSE"),
    .CLKIN_PERIOD          (125.0),
    .CLKFX_MD_MAX          (0.000))
   dcm_clkgen_inst
    // Input clock
   (.CLKIN                 (clk_8),
    // Output clocks
    .CLKFX                 (clkgen),
    // Ports for dynamic reconfiguration
    .PROGCLK               (clk_ref),
    .PROGDATA              (prog_data[0]),
    .PROGEN                (prog_en[0]),
    .PROGDONE              (prog_done),
    // Other control and status signals
    .FREEZEDCM             (1'b0),
    .LOCKED                (locked_dcm),
    .STATUS                (),
    .RST                   (reset)
);

// input freq to pll (28 or generated from 8)
wire clkpllin;
BUFGMUX clk_in_mux(.I0(clk_ref), .I1(clkgen), .O(clkpllin), .S(vdac2_sel));

// pll resetter
wire pll_rst;
pll_reset pll_reset(
	.clk(clk_ref),
	.i_reset((vdac2_sel) ? (~locked_dcm || reset) : (hdmi_reset || reset)),
	.o_reset(pll_rst)
);
assign o_reset = pll_rst;

// pll to produce x5 clock
wire clk0, clkfx, clkfx180, clkdv, clkfbout, lockedx5;

DCM_SP
  #(.CLKDV_DIVIDE          (2.000),
    .CLKFX_DIVIDE          (1),
    .CLKFX_MULTIPLY        (5),
    .CLKIN_DIVIDE_BY_2     ("FALSE"),
    .CLKIN_PERIOD          (13.000),
    .CLKOUT_PHASE_SHIFT    ("NONE"),
    .CLK_FEEDBACK          ("1X"),
    .DESKEW_ADJUST         ("SYSTEM_SYNCHRONOUS"),
    .PHASE_SHIFT           (0),
    .STARTUP_WAIT          ("FALSE"))
  dcm_sp_inst
    // Input clock
   (.CLKIN                 (clkpllin),
    .CLKFB                 (clkfbout),
    // Output clocks
    .CLK0                  (clk0),
    .CLK90                 (),
    .CLK180                (),
    .CLK270                (),
    .CLK2X                 (),
    .CLK2X180              (),
    .CLKFX                 (clkfx),
    .CLKFX180              (clkfx180),
    .CLKDV                 (clkdv),
    // Ports for dynamic phase shift
    .PSCLK                 (1'b0),
    .PSEN                  (1'b0),
    .PSINCDEC              (1'b0),
    .PSDONE                (),
    // Other control and status signals
    .LOCKED                (lockedx5),
    .STATUS                (),
    .RST                   (pll_rst),
    .DSSEN                 (1'b0));

// feedback buf
BUFG clkf_buf(.O (clkfbout), .I (clk0));

// output bufs
BUFG clkout1_buf (.O(clk_hdmi), .I(clkfx));
BUFG clkout2_buf (.O(clk_hdmi_n), .I(clkfx180));
BUFG clkout3_buf (.O(clk_pix), .I(clk0));
BUFG clkout4_buf (.O(clk_pix2), .I(clkdv));
assign locked = lockedx5;

endmodule
