//============================================================================
//  Audio compressor (signed samples)
// 
//  Copyright (C) 2018 Sorgelig
//  Converted to verilog (c) 2025 Andy Karpov
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//
//  You should have received a copy of the GNU General Public License along
//  with this program; if not, write to the Free Software Foundation, Inc.,
//  51 Franklin Street, Fifth Floor, Boston, MA 02110-1301 USA.
//============================================================================

module compressor
(
	input wire clk,
	input wire [11:0] in1, in2,
	output reg [15:0] out1, out2
);

always @(posedge clk) out1 <= {in1[11], in1[11] ? ~tbl[~in1[10:0]] : tbl[in1[10:0]]};
always @(posedge clk) out2 <= {in2[11], in2[11] ? ~tbl[~in2[10:0]] : tbl[in2[10:0]]};

reg[14:0] tbl[0:2047];
initial begin 
	tbl[0] = 15'h0000;
	tbl[1] = 15'h0019;
	tbl[2] = 15'h0032;
	tbl[3] = 15'h004B;
	tbl[4] = 15'h0064;
	tbl[5] = 15'h007D;
	tbl[6] = 15'h0096;
	tbl[7] = 15'h00B0;
	tbl[8] = 15'h00C9;
	tbl[9] = 15'h00E2;
	tbl[10] = 15'h00FB;
	tbl[11] = 15'h0114;
	tbl[12] = 15'h012D;
	tbl[13] = 15'h0146;
	tbl[14] = 15'h0160;
	tbl[15] = 15'h0179;
	tbl[16] = 15'h0192;
	tbl[17] = 15'h01AB;
	tbl[18] = 15'h01C4;
	tbl[19] = 15'h01DD;
	tbl[20] = 15'h01F6;
	tbl[21] = 15'h0210;
	tbl[22] = 15'h0229;
	tbl[23] = 15'h0242;
	tbl[24] = 15'h025B;
	tbl[25] = 15'h0274;
	tbl[26] = 15'h028D;
	tbl[27] = 15'h02A6;
	tbl[28] = 15'h02BF;
	tbl[29] = 15'h02D9;
	tbl[30] = 15'h02F2;
	tbl[31] = 15'h030B;
	tbl[32] = 15'h0324;
	tbl[33] = 15'h033D;
	tbl[34] = 15'h0356;
	tbl[35] = 15'h036F;
	tbl[36] = 15'h0389;
	tbl[37] = 15'h03A2;
	tbl[38] = 15'h03BB;
	tbl[39] = 15'h03D4;
	tbl[40] = 15'h03ED;
	tbl[41] = 15'h0406;
	tbl[42] = 15'h041F;
	tbl[43] = 15'h0439;
	tbl[44] = 15'h0452;
	tbl[45] = 15'h046B;
	tbl[46] = 15'h0484;
	tbl[47] = 15'h049D;
	tbl[48] = 15'h04B6;
	tbl[49] = 15'h04CF;
	tbl[50] = 15'h04E8;
	tbl[51] = 15'h0502;
	tbl[52] = 15'h051B;
	tbl[53] = 15'h0534;
	tbl[54] = 15'h054D;
	tbl[55] = 15'h0566;
	tbl[56] = 15'h057F;
	tbl[57] = 15'h0598;
	tbl[58] = 15'h05B1;
	tbl[59] = 15'h05CB;
	tbl[60] = 15'h05E4;
	tbl[61] = 15'h05FD;
	tbl[62] = 15'h0616;
	tbl[63] = 15'h062F;
	tbl[64] = 15'h0648;
	tbl[65] = 15'h0661;
	tbl[66] = 15'h067A;
	tbl[67] = 15'h0693;
	tbl[68] = 15'h06AD;
	tbl[69] = 15'h06C6;
	tbl[70] = 15'h06DF;
	tbl[71] = 15'h06F8;
	tbl[72] = 15'h0711;
	tbl[73] = 15'h072A;
	tbl[74] = 15'h0743;
	tbl[75] = 15'h075C;
	tbl[76] = 15'h0775;
	tbl[77] = 15'h078E;
	tbl[78] = 15'h07A8;
	tbl[79] = 15'h07C1;
	tbl[80] = 15'h07DA;
	tbl[81] = 15'h07F3;
	tbl[82] = 15'h080C;
	tbl[83] = 15'h0825;
	tbl[84] = 15'h083E;
	tbl[85] = 15'h0857;
	tbl[86] = 15'h0870;
	tbl[87] = 15'h0889;
	tbl[88] = 15'h08A3;
	tbl[89] = 15'h08BC;
	tbl[90] = 15'h08D5;
	tbl[91] = 15'h08EE;
	tbl[92] = 15'h0907;
	tbl[93] = 15'h0920;
	tbl[94] = 15'h0939;
	tbl[95] = 15'h0952;
	tbl[96] = 15'h096B;
	tbl[97] = 15'h0984;
	tbl[98] = 15'h099D;
	tbl[99] = 15'h09B6;
	tbl[100] = 15'h09CF;
	tbl[101] = 15'h09E9;
	tbl[102] = 15'h0A02;
	tbl[103] = 15'h0A1B;
	tbl[104] = 15'h0A34;
	tbl[105] = 15'h0A4D;
	tbl[106] = 15'h0A66;
	tbl[107] = 15'h0A7F;
	tbl[108] = 15'h0A98;
	tbl[109] = 15'h0AB1;
	tbl[110] = 15'h0ACA;
	tbl[111] = 15'h0AE3;
	tbl[112] = 15'h0AFC;
	tbl[113] = 15'h0B15;
	tbl[114] = 15'h0B2E;
	tbl[115] = 15'h0B47;
	tbl[116] = 15'h0B60;
	tbl[117] = 15'h0B79;
	tbl[118] = 15'h0B92;
	tbl[119] = 15'h0BAC;
	tbl[120] = 15'h0BC5;
	tbl[121] = 15'h0BDE;
	tbl[122] = 15'h0BF7;
	tbl[123] = 15'h0C10;
	tbl[124] = 15'h0C29;
	tbl[125] = 15'h0C42;
	tbl[126] = 15'h0C5B;
	tbl[127] = 15'h0C74;
	tbl[128] = 15'h0C8D;
	tbl[129] = 15'h0CA6;
	tbl[130] = 15'h0CBF;
	tbl[131] = 15'h0CD8;
	tbl[132] = 15'h0CF1;
	tbl[133] = 15'h0D0A;
	tbl[134] = 15'h0D23;
	tbl[135] = 15'h0D3C;
	tbl[136] = 15'h0D55;
	tbl[137] = 15'h0D6E;
	tbl[138] = 15'h0D87;
	tbl[139] = 15'h0DA0;
	tbl[140] = 15'h0DB9;
	tbl[141] = 15'h0DD2;
	tbl[142] = 15'h0DEB;
	tbl[143] = 15'h0E04;
	tbl[144] = 15'h0E1D;
	tbl[145] = 15'h0E36;
	tbl[146] = 15'h0E4F;
	tbl[147] = 15'h0E68;
	tbl[148] = 15'h0E81;
	tbl[149] = 15'h0E9A;
	tbl[150] = 15'h0EB3;
	tbl[151] = 15'h0ECC;
	tbl[152] = 15'h0EE5;
	tbl[153] = 15'h0EFE;
	tbl[154] = 15'h0F17;
	tbl[155] = 15'h0F30;
	tbl[156] = 15'h0F49;
	tbl[157] = 15'h0F62;
	tbl[158] = 15'h0F7B;
	tbl[159] = 15'h0F94;
	tbl[160] = 15'h0FAC;
	tbl[161] = 15'h0FC5;
	tbl[162] = 15'h0FDE;
	tbl[163] = 15'h0FF7;
	tbl[164] = 15'h1010;
	tbl[165] = 15'h1029;
	tbl[166] = 15'h1042;
	tbl[167] = 15'h105B;
	tbl[168] = 15'h1074;
	tbl[169] = 15'h108D;
	tbl[170] = 15'h10A6;
	tbl[171] = 15'h10BF;
	tbl[172] = 15'h10D8;
	tbl[173] = 15'h10F1;
	tbl[174] = 15'h110A;
	tbl[175] = 15'h1123;
	tbl[176] = 15'h113B;
	tbl[177] = 15'h1154;
	tbl[178] = 15'h116D;
	tbl[179] = 15'h1186;
	tbl[180] = 15'h119F;
	tbl[181] = 15'h11B8;
	tbl[182] = 15'h11D1;
	tbl[183] = 15'h11EA;
	tbl[184] = 15'h1203;
	tbl[185] = 15'h121C;
	tbl[186] = 15'h1234;
	tbl[187] = 15'h124D;
	tbl[188] = 15'h1266;
	tbl[189] = 15'h127F;
	tbl[190] = 15'h1298;
	tbl[191] = 15'h12B1;
	tbl[192] = 15'h12CA;
	tbl[193] = 15'h12E3;
	tbl[194] = 15'h12FB;
	tbl[195] = 15'h1314;
	tbl[196] = 15'h132D;
	tbl[197] = 15'h1346;
	tbl[198] = 15'h135F;
	tbl[199] = 15'h1378;
	tbl[200] = 15'h1391;
	tbl[201] = 15'h13A9;
	tbl[202] = 15'h13C2;
	tbl[203] = 15'h13DB;
	tbl[204] = 15'h13F4;
	tbl[205] = 15'h140D;
	tbl[206] = 15'h1426;
	tbl[207] = 15'h143E;
	tbl[208] = 15'h1457;
	tbl[209] = 15'h1470;
	tbl[210] = 15'h1489;
	tbl[211] = 15'h14A2;
	tbl[212] = 15'h14BB;
	tbl[213] = 15'h14D3;
	tbl[214] = 15'h14EC;
	tbl[215] = 15'h1505;
	tbl[216] = 15'h151E;
	tbl[217] = 15'h1537;
	tbl[218] = 15'h154F;
	tbl[219] = 15'h1568;
	tbl[220] = 15'h1581;
	tbl[221] = 15'h159A;
	tbl[222] = 15'h15B3;
	tbl[223] = 15'h15CB;
	tbl[224] = 15'h15E4;
	tbl[225] = 15'h15FD;
	tbl[226] = 15'h1616;
	tbl[227] = 15'h162E;
	tbl[228] = 15'h1647;
	tbl[229] = 15'h1660;
	tbl[230] = 15'h1679;
	tbl[231] = 15'h1691;
	tbl[232] = 15'h16AA;
	tbl[233] = 15'h16C3;
	tbl[234] = 15'h16DC;
	tbl[235] = 15'h16F4;
	tbl[236] = 15'h170D;
	tbl[237] = 15'h1726;
	tbl[238] = 15'h173F;
	tbl[239] = 15'h1757;
	tbl[240] = 15'h1770;
	tbl[241] = 15'h1789;
	tbl[242] = 15'h17A1;
	tbl[243] = 15'h17BA;
	tbl[244] = 15'h17D3;
	tbl[245] = 15'h17EC;
	tbl[246] = 15'h1804;
	tbl[247] = 15'h181D;
	tbl[248] = 15'h1836;
	tbl[249] = 15'h184E;
	tbl[250] = 15'h1867;
	tbl[251] = 15'h1880;
	tbl[252] = 15'h1898;
	tbl[253] = 15'h18B1;
	tbl[254] = 15'h18CA;
	tbl[255] = 15'h18E2;
	tbl[256] = 15'h18FB;
	tbl[257] = 15'h1914;
	tbl[258] = 15'h192C;
	tbl[259] = 15'h1945;
	tbl[260] = 15'h195E;
	tbl[261] = 15'h1976;
	tbl[262] = 15'h198F;
	tbl[263] = 15'h19A8;
	tbl[264] = 15'h19C0;
	tbl[265] = 15'h19D9;
	tbl[266] = 15'h19F2;
	tbl[267] = 15'h1A0A;
	tbl[268] = 15'h1A23;
	tbl[269] = 15'h1A3B;
	tbl[270] = 15'h1A54;
	tbl[271] = 15'h1A6D;
	tbl[272] = 15'h1A85;
	tbl[273] = 15'h1A9E;
	tbl[274] = 15'h1AB6;
	tbl[275] = 15'h1ACF;
	tbl[276] = 15'h1AE8;
	tbl[277] = 15'h1B00;
	tbl[278] = 15'h1B19;
	tbl[279] = 15'h1B31;
	tbl[280] = 15'h1B4A;
	tbl[281] = 15'h1B62;
	tbl[282] = 15'h1B7B;
	tbl[283] = 15'h1B94;
	tbl[284] = 15'h1BAC;
	tbl[285] = 15'h1BC5;
	tbl[286] = 15'h1BDD;
	tbl[287] = 15'h1BF6;
	tbl[288] = 15'h1C0E;
	tbl[289] = 15'h1C27;
	tbl[290] = 15'h1C3F;
	tbl[291] = 15'h1C58;
	tbl[292] = 15'h1C70;
	tbl[293] = 15'h1C89;
	tbl[294] = 15'h1CA1;
	tbl[295] = 15'h1CBA;
	tbl[296] = 15'h1CD2;
	tbl[297] = 15'h1CEB;
	tbl[298] = 15'h1D03;
	tbl[299] = 15'h1D1C;
	tbl[300] = 15'h1D34;
	tbl[301] = 15'h1D4D;
	tbl[302] = 15'h1D65;
	tbl[303] = 15'h1D7E;
	tbl[304] = 15'h1D96;
	tbl[305] = 15'h1DAF;
	tbl[306] = 15'h1DC7;
	tbl[307] = 15'h1DE0;
	tbl[308] = 15'h1DF8;
	tbl[309] = 15'h1E10;
	tbl[310] = 15'h1E29;
	tbl[311] = 15'h1E41;
	tbl[312] = 15'h1E5A;
	tbl[313] = 15'h1E72;
	tbl[314] = 15'h1E8B;
	tbl[315] = 15'h1EA3;
	tbl[316] = 15'h1EBB;
	tbl[317] = 15'h1ED4;
	tbl[318] = 15'h1EEC;
	tbl[319] = 15'h1F05;
	tbl[320] = 15'h1F1D;
	tbl[321] = 15'h1F35;
	tbl[322] = 15'h1F4E;
	tbl[323] = 15'h1F66;
	tbl[324] = 15'h1F7F;
	tbl[325] = 15'h1F97;
	tbl[326] = 15'h1FAF;
	tbl[327] = 15'h1FC8;
	tbl[328] = 15'h1FE0;
	tbl[329] = 15'h1FF8;
	tbl[330] = 15'h2011;
	tbl[331] = 15'h2029;
	tbl[332] = 15'h2041;
	tbl[333] = 15'h205A;
	tbl[334] = 15'h2072;
	tbl[335] = 15'h208A;
	tbl[336] = 15'h20A3;
	tbl[337] = 15'h20BB;
	tbl[338] = 15'h20D3;
	tbl[339] = 15'h20EC;
	tbl[340] = 15'h2104;
	tbl[341] = 15'h211C;
	tbl[342] = 15'h2134;
	tbl[343] = 15'h214D;
	tbl[344] = 15'h2165;
	tbl[345] = 15'h217D;
	tbl[346] = 15'h2196;
	tbl[347] = 15'h21AE;
	tbl[348] = 15'h21C6;
	tbl[349] = 15'h21DE;
	tbl[350] = 15'h21F7;
	tbl[351] = 15'h220F;
	tbl[352] = 15'h2227;
	tbl[353] = 15'h223F;
	tbl[354] = 15'h2257;
	tbl[355] = 15'h2270;
	tbl[356] = 15'h2288;
	tbl[357] = 15'h22A0;
	tbl[358] = 15'h22B8;
	tbl[359] = 15'h22D1;
	tbl[360] = 15'h22E9;
	tbl[361] = 15'h2301;
	tbl[362] = 15'h2319;
	tbl[363] = 15'h2331;
	tbl[364] = 15'h2349;
	tbl[365] = 15'h2362;
	tbl[366] = 15'h237A;
	tbl[367] = 15'h2392;
	tbl[368] = 15'h23AA;
	tbl[369] = 15'h23C2;
	tbl[370] = 15'h23DA;
	tbl[371] = 15'h23F3;
	tbl[372] = 15'h240B;
	tbl[373] = 15'h2423;
	tbl[374] = 15'h243B;
	tbl[375] = 15'h2453;
	tbl[376] = 15'h246B;
	tbl[377] = 15'h2483;
	tbl[378] = 15'h249B;
	tbl[379] = 15'h24B3;
	tbl[380] = 15'h24CB;
	tbl[381] = 15'h24E4;
	tbl[382] = 15'h24FC;
	tbl[383] = 15'h2514;
	tbl[384] = 15'h252C;
	tbl[385] = 15'h2544;
	tbl[386] = 15'h255C;
	tbl[387] = 15'h2574;
	tbl[388] = 15'h258C;
	tbl[389] = 15'h25A4;
	tbl[390] = 15'h25BC;
	tbl[391] = 15'h25D4;
	tbl[392] = 15'h25EC;
	tbl[393] = 15'h2604;
	tbl[394] = 15'h261C;
	tbl[395] = 15'h2634;
	tbl[396] = 15'h264C;
	tbl[397] = 15'h2664;
	tbl[398] = 15'h267C;
	tbl[399] = 15'h2694;
	tbl[400] = 15'h26AC;
	tbl[401] = 15'h26C4;
	tbl[402] = 15'h26DC;
	tbl[403] = 15'h26F4;
	tbl[404] = 15'h270C;
	tbl[405] = 15'h2724;
	tbl[406] = 15'h273C;
	tbl[407] = 15'h2754;
	tbl[408] = 15'h276C;
	tbl[409] = 15'h2783;
	tbl[410] = 15'h279B;
	tbl[411] = 15'h27B3;
	tbl[412] = 15'h27CB;
	tbl[413] = 15'h27E3;
	tbl[414] = 15'h27FB;
	tbl[415] = 15'h2813;
	tbl[416] = 15'h282B;
	tbl[417] = 15'h2843;
	tbl[418] = 15'h285A;
	tbl[419] = 15'h2872;
	tbl[420] = 15'h288A;
	tbl[421] = 15'h28A2;
	tbl[422] = 15'h28BA;
	tbl[423] = 15'h28D2;
	tbl[424] = 15'h28EA;
	tbl[425] = 15'h2901;
	tbl[426] = 15'h2919;
	tbl[427] = 15'h2931;
	tbl[428] = 15'h2949;
	tbl[429] = 15'h2961;
	tbl[430] = 15'h2978;
	tbl[431] = 15'h2990;
	tbl[432] = 15'h29A8;
	tbl[433] = 15'h29C0;
	tbl[434] = 15'h29D7;
	tbl[435] = 15'h29EF;
	tbl[436] = 15'h2A07;
	tbl[437] = 15'h2A1F;
	tbl[438] = 15'h2A36;
	tbl[439] = 15'h2A4E;
	tbl[440] = 15'h2A66;
	tbl[441] = 15'h2A7E;
	tbl[442] = 15'h2A95;
	tbl[443] = 15'h2AAD;
	tbl[444] = 15'h2AC5;
	tbl[445] = 15'h2ADC;
	tbl[446] = 15'h2AF4;
	tbl[447] = 15'h2B0C;
	tbl[448] = 15'h2B24;
	tbl[449] = 15'h2B3B;
	tbl[450] = 15'h2B53;
	tbl[451] = 15'h2B6B;
	tbl[452] = 15'h2B82;
	tbl[453] = 15'h2B9A;
	tbl[454] = 15'h2BB1;
	tbl[455] = 15'h2BC9;
	tbl[456] = 15'h2BE1;
	tbl[457] = 15'h2BF8;
	tbl[458] = 15'h2C10;
	tbl[459] = 15'h2C28;
	tbl[460] = 15'h2C3F;
	tbl[461] = 15'h2C57;
	tbl[462] = 15'h2C6E;
	tbl[463] = 15'h2C86;
	tbl[464] = 15'h2C9D;
	tbl[465] = 15'h2CB5;
	tbl[466] = 15'h2CCD;
	tbl[467] = 15'h2CE4;
	tbl[468] = 15'h2CFC;
	tbl[469] = 15'h2D13;
	tbl[470] = 15'h2D2B;
	tbl[471] = 15'h2D42;
	tbl[472] = 15'h2D5A;
	tbl[473] = 15'h2D71;
	tbl[474] = 15'h2D89;
	tbl[475] = 15'h2DA0;
	tbl[476] = 15'h2DB8;
	tbl[477] = 15'h2DCF;
	tbl[478] = 15'h2DE7;
	tbl[479] = 15'h2DFE;
	tbl[480] = 15'h2E16;
	tbl[481] = 15'h2E2D;
	tbl[482] = 15'h2E45;
	tbl[483] = 15'h2E5C;
	tbl[484] = 15'h2E73;
	tbl[485] = 15'h2E8B;
	tbl[486] = 15'h2EA2;
	tbl[487] = 15'h2EBA;
	tbl[488] = 15'h2ED1;
	tbl[489] = 15'h2EE9;
	tbl[490] = 15'h2F00;
	tbl[491] = 15'h2F17;
	tbl[492] = 15'h2F2F;
	tbl[493] = 15'h2F46;
	tbl[494] = 15'h2F5D;
	tbl[495] = 15'h2F75;
	tbl[496] = 15'h2F8C;
	tbl[497] = 15'h2FA3;
	tbl[498] = 15'h2FBB;
	tbl[499] = 15'h2FD2;
	tbl[500] = 15'h2FE9;
	tbl[501] = 15'h3001;
	tbl[502] = 15'h3018;
	tbl[503] = 15'h302F;
	tbl[504] = 15'h3047;
	tbl[505] = 15'h305E;
	tbl[506] = 15'h3075;
	tbl[507] = 15'h308C;
	tbl[508] = 15'h30A4;
	tbl[509] = 15'h30BB;
	tbl[510] = 15'h30D2;
	tbl[511] = 15'h30E9;
	tbl[512] = 15'h3101;
	tbl[513] = 15'h3118;
	tbl[514] = 15'h312F;
	tbl[515] = 15'h3146;
	tbl[516] = 15'h315E;
	tbl[517] = 15'h3175;
	tbl[518] = 15'h318C;
	tbl[519] = 15'h31A3;
	tbl[520] = 15'h31BA;
	tbl[521] = 15'h31D1;
	tbl[522] = 15'h31E9;
	tbl[523] = 15'h3200;
	tbl[524] = 15'h3217;
	tbl[525] = 15'h322E;
	tbl[526] = 15'h3245;
	tbl[527] = 15'h325C;
	tbl[528] = 15'h3273;
	tbl[529] = 15'h328A;
	tbl[530] = 15'h32A2;
	tbl[531] = 15'h32B9;
	tbl[532] = 15'h32D0;
	tbl[533] = 15'h32E7;
	tbl[534] = 15'h32FE;
	tbl[535] = 15'h3315;
	tbl[536] = 15'h332C;
	tbl[537] = 15'h3343;
	tbl[538] = 15'h335A;
	tbl[539] = 15'h3371;
	tbl[540] = 15'h3388;
	tbl[541] = 15'h339F;
	tbl[542] = 15'h33B6;
	tbl[543] = 15'h33CD;
	tbl[544] = 15'h33E4;
	tbl[545] = 15'h33FB;
	tbl[546] = 15'h3412;
	tbl[547] = 15'h3429;
	tbl[548] = 15'h3440;
	tbl[549] = 15'h3457;
	tbl[550] = 15'h346E;
	tbl[551] = 15'h3485;
	tbl[552] = 15'h349C;
	tbl[553] = 15'h34B3;
	tbl[554] = 15'h34CA;
	tbl[555] = 15'h34E1;
	tbl[556] = 15'h34F7;
	tbl[557] = 15'h350E;
	tbl[558] = 15'h3525;
	tbl[559] = 15'h353C;
	tbl[560] = 15'h3553;
	tbl[561] = 15'h356A;
	tbl[562] = 15'h3581;
	tbl[563] = 15'h3597;
	tbl[564] = 15'h35AE;
	tbl[565] = 15'h35C5;
	tbl[566] = 15'h35DC;
	tbl[567] = 15'h35F3;
	tbl[568] = 15'h360A;
	tbl[569] = 15'h3620;
	tbl[570] = 15'h3637;
	tbl[571] = 15'h364E;
	tbl[572] = 15'h3665;
	tbl[573] = 15'h367B;
	tbl[574] = 15'h3692;
	tbl[575] = 15'h36A9;
	tbl[576] = 15'h36C0;
	tbl[577] = 15'h36D6;
	tbl[578] = 15'h36ED;
	tbl[579] = 15'h3704;
	tbl[580] = 15'h371A;
	tbl[581] = 15'h3731;
	tbl[582] = 15'h3748;
	tbl[583] = 15'h375E;
	tbl[584] = 15'h3775;
	tbl[585] = 15'h378C;
	tbl[586] = 15'h37A2;
	tbl[587] = 15'h37B9;
	tbl[588] = 15'h37D0;
	tbl[589] = 15'h37E6;
	tbl[590] = 15'h37FD;
	tbl[591] = 15'h3814;
	tbl[592] = 15'h382A;
	tbl[593] = 15'h3841;
	tbl[594] = 15'h3857;
	tbl[595] = 15'h386E;
	tbl[596] = 15'h3884;
	tbl[597] = 15'h389B;
	tbl[598] = 15'h38B2;
	tbl[599] = 15'h38C8;
	tbl[600] = 15'h38DF;
	tbl[601] = 15'h38F5;
	tbl[602] = 15'h390C;
	tbl[603] = 15'h3922;
	tbl[604] = 15'h3939;
	tbl[605] = 15'h394F;
	tbl[606] = 15'h3966;
	tbl[607] = 15'h397C;
	tbl[608] = 15'h3993;
	tbl[609] = 15'h39A9;
	tbl[610] = 15'h39BF;
	tbl[611] = 15'h39D6;
	tbl[612] = 15'h39EC;
	tbl[613] = 15'h3A03;
	tbl[614] = 15'h3A19;
	tbl[615] = 15'h3A30;
	tbl[616] = 15'h3A46;
	tbl[617] = 15'h3A5C;
	tbl[618] = 15'h3A73;
	tbl[619] = 15'h3A89;
	tbl[620] = 15'h3A9F;
	tbl[621] = 15'h3AB6;
	tbl[622] = 15'h3ACC;
	tbl[623] = 15'h3AE2;
	tbl[624] = 15'h3AF9;
	tbl[625] = 15'h3B0F;
	tbl[626] = 15'h3B25;
	tbl[627] = 15'h3B3C;
	tbl[628] = 15'h3B52;
	tbl[629] = 15'h3B68;
	tbl[630] = 15'h3B7F;
	tbl[631] = 15'h3B95;
	tbl[632] = 15'h3BAB;
	tbl[633] = 15'h3BC1;
	tbl[634] = 15'h3BD7;
	tbl[635] = 15'h3BEE;
	tbl[636] = 15'h3C04;
	tbl[637] = 15'h3C1A;
	tbl[638] = 15'h3C30;
	tbl[639] = 15'h3C47;
	tbl[640] = 15'h3C5D;
	tbl[641] = 15'h3C73;
	tbl[642] = 15'h3C89;
	tbl[643] = 15'h3C9F;
	tbl[644] = 15'h3CB5;
	tbl[645] = 15'h3CCB;
	tbl[646] = 15'h3CE2;
	tbl[647] = 15'h3CF8;
	tbl[648] = 15'h3D0E;
	tbl[649] = 15'h3D24;
	tbl[650] = 15'h3D3A;
	tbl[651] = 15'h3D50;
	tbl[652] = 15'h3D66;
	tbl[653] = 15'h3D7C;
	tbl[654] = 15'h3D92;
	tbl[655] = 15'h3DA8;
	tbl[656] = 15'h3DBE;
	tbl[657] = 15'h3DD4;
	tbl[658] = 15'h3DEA;
	tbl[659] = 15'h3E00;
	tbl[660] = 15'h3E16;
	tbl[661] = 15'h3E2C;
	tbl[662] = 15'h3E42;
	tbl[663] = 15'h3E58;
	tbl[664] = 15'h3E6E;
	tbl[665] = 15'h3E84;
	tbl[666] = 15'h3E9A;
	tbl[667] = 15'h3EB0;
	tbl[668] = 15'h3EC6;
	tbl[669] = 15'h3EDC;
	tbl[670] = 15'h3EF2;
	tbl[671] = 15'h3F08;
	tbl[672] = 15'h3F1D;
	tbl[673] = 15'h3F33;
	tbl[674] = 15'h3F49;
	tbl[675] = 15'h3F5F;
	tbl[676] = 15'h3F75;
	tbl[677] = 15'h3F8B;
	tbl[678] = 15'h3FA1;
	tbl[679] = 15'h3FB6;
	tbl[680] = 15'h3FCC;
	tbl[681] = 15'h3FE2;
	tbl[682] = 15'h3FF8;
	tbl[683] = 15'h400E;
	tbl[684] = 15'h4023;
	tbl[685] = 15'h4039;
	tbl[686] = 15'h404F;
	tbl[687] = 15'h4065;
	tbl[688] = 15'h407A;
	tbl[689] = 15'h4090;
	tbl[690] = 15'h40A6;
	tbl[691] = 15'h40BB;
	tbl[692] = 15'h40D1;
	tbl[693] = 15'h40E7;
	tbl[694] = 15'h40FC;
	tbl[695] = 15'h4112;
	tbl[696] = 15'h4128;
	tbl[697] = 15'h413D;
	tbl[698] = 15'h4153;
	tbl[699] = 15'h4169;
	tbl[700] = 15'h417E;
	tbl[701] = 15'h4194;
	tbl[702] = 15'h41A9;
	tbl[703] = 15'h41BF;
	tbl[704] = 15'h41D5;
	tbl[705] = 15'h41EA;
	tbl[706] = 15'h4200;
	tbl[707] = 15'h4215;
	tbl[708] = 15'h422B;
	tbl[709] = 15'h4240;
	tbl[710] = 15'h4256;
	tbl[711] = 15'h426B;
	tbl[712] = 15'h4281;
	tbl[713] = 15'h4296;
	tbl[714] = 15'h42AC;
	tbl[715] = 15'h42C1;
	tbl[716] = 15'h42D7;
	tbl[717] = 15'h42EC;
	tbl[718] = 15'h4301;
	tbl[719] = 15'h4317;
	tbl[720] = 15'h432C;
	tbl[721] = 15'h4342;
	tbl[722] = 15'h4357;
	tbl[723] = 15'h436C;
	tbl[724] = 15'h4382;
	tbl[725] = 15'h4397;
	tbl[726] = 15'h43AC;
	tbl[727] = 15'h43C2;
	tbl[728] = 15'h43D7;
	tbl[729] = 15'h43EC;
	tbl[730] = 15'h4402;
	tbl[731] = 15'h4417;
	tbl[732] = 15'h442C;
	tbl[733] = 15'h4442;
	tbl[734] = 15'h4457;
	tbl[735] = 15'h446C;
	tbl[736] = 15'h4481;
	tbl[737] = 15'h4497;
	tbl[738] = 15'h44AC;
	tbl[739] = 15'h44C1;
	tbl[740] = 15'h44D6;
	tbl[741] = 15'h44EB;
	tbl[742] = 15'h4501;
	tbl[743] = 15'h4516;
	tbl[744] = 15'h452B;
	tbl[745] = 15'h4540;
	tbl[746] = 15'h4555;
	tbl[747] = 15'h456A;
	tbl[748] = 15'h4580;
	tbl[749] = 15'h4595;
	tbl[750] = 15'h45AA;
	tbl[751] = 15'h45BF;
	tbl[752] = 15'h45D4;
	tbl[753] = 15'h45E9;
	tbl[754] = 15'h45FE;
	tbl[755] = 15'h4613;
	tbl[756] = 15'h4628;
	tbl[757] = 15'h463D;
	tbl[758] = 15'h4652;
	tbl[759] = 15'h4667;
	tbl[760] = 15'h467C;
	tbl[761] = 15'h4691;
	tbl[762] = 15'h46A6;
	tbl[763] = 15'h46BB;
	tbl[764] = 15'h46D0;
	tbl[765] = 15'h46E5;
	tbl[766] = 15'h46FA;
	tbl[767] = 15'h470F;
	tbl[768] = 15'h4724;
	tbl[769] = 15'h4739;
	tbl[770] = 15'h474D;
	tbl[771] = 15'h4762;
	tbl[772] = 15'h4777;
	tbl[773] = 15'h478C;
	tbl[774] = 15'h47A1;
	tbl[775] = 15'h47B6;
	tbl[776] = 15'h47CB;
	tbl[777] = 15'h47DF;
	tbl[778] = 15'h47F4;
	tbl[779] = 15'h4809;
	tbl[780] = 15'h481E;
	tbl[781] = 15'h4833;
	tbl[782] = 15'h4847;
	tbl[783] = 15'h485C;
	tbl[784] = 15'h4871;
	tbl[785] = 15'h4885;
	tbl[786] = 15'h489A;
	tbl[787] = 15'h48AF;
	tbl[788] = 15'h48C4;
	tbl[789] = 15'h48D8;
	tbl[790] = 15'h48ED;
	tbl[791] = 15'h4902;
	tbl[792] = 15'h4916;
	tbl[793] = 15'h492B;
	tbl[794] = 15'h4940;
	tbl[795] = 15'h4954;
	tbl[796] = 15'h4969;
	tbl[797] = 15'h497D;
	tbl[798] = 15'h4992;
	tbl[799] = 15'h49A6;
	tbl[800] = 15'h49BB;
	tbl[801] = 15'h49D0;
	tbl[802] = 15'h49E4;
	tbl[803] = 15'h49F9;
	tbl[804] = 15'h4A0D;
	tbl[805] = 15'h4A22;
	tbl[806] = 15'h4A36;
	tbl[807] = 15'h4A4B;
	tbl[808] = 15'h4A5F;
	tbl[809] = 15'h4A74;
	tbl[810] = 15'h4A88;
	tbl[811] = 15'h4A9C;
	tbl[812] = 15'h4AB1;
	tbl[813] = 15'h4AC5;
	tbl[814] = 15'h4ADA;
	tbl[815] = 15'h4AEE;
	tbl[816] = 15'h4B02;
	tbl[817] = 15'h4B17;
	tbl[818] = 15'h4B2B;
	tbl[819] = 15'h4B40;
	tbl[820] = 15'h4B54;
	tbl[821] = 15'h4B68;
	tbl[822] = 15'h4B7C;
	tbl[823] = 15'h4B91;
	tbl[824] = 15'h4BA5;
	tbl[825] = 15'h4BB9;
	tbl[826] = 15'h4BCE;
	tbl[827] = 15'h4BE2;
	tbl[828] = 15'h4BF6;
	tbl[829] = 15'h4C0A;
	tbl[830] = 15'h4C1F;
	tbl[831] = 15'h4C33;
	tbl[832] = 15'h4C47;
	tbl[833] = 15'h4C5B;
	tbl[834] = 15'h4C6F;
	tbl[835] = 15'h4C84;
	tbl[836] = 15'h4C98;
	tbl[837] = 15'h4CAC;
	tbl[838] = 15'h4CC0;
	tbl[839] = 15'h4CD4;
	tbl[840] = 15'h4CE8;
	tbl[841] = 15'h4CFC;
	tbl[842] = 15'h4D10;
	tbl[843] = 15'h4D24;
	tbl[844] = 15'h4D38;
	tbl[845] = 15'h4D4C;
	tbl[846] = 15'h4D61;
	tbl[847] = 15'h4D75;
	tbl[848] = 15'h4D89;
	tbl[849] = 15'h4D9D;
	tbl[850] = 15'h4DB1;
	tbl[851] = 15'h4DC5;
	tbl[852] = 15'h4DD8;
	tbl[853] = 15'h4DEC;
	tbl[854] = 15'h4E00;
	tbl[855] = 15'h4E14;
	tbl[856] = 15'h4E28;
	tbl[857] = 15'h4E3C;
	tbl[858] = 15'h4E50;
	tbl[859] = 15'h4E64;
	tbl[860] = 15'h4E78;
	tbl[861] = 15'h4E8C;
	tbl[862] = 15'h4E9F;
	tbl[863] = 15'h4EB3;
	tbl[864] = 15'h4EC7;
	tbl[865] = 15'h4EDB;
	tbl[866] = 15'h4EEF;
	tbl[867] = 15'h4F03;
	tbl[868] = 15'h4F16;
	tbl[869] = 15'h4F2A;
	tbl[870] = 15'h4F3E;
	tbl[871] = 15'h4F52;
	tbl[872] = 15'h4F65;
	tbl[873] = 15'h4F79;
	tbl[874] = 15'h4F8D;
	tbl[875] = 15'h4FA0;
	tbl[876] = 15'h4FB4;
	tbl[877] = 15'h4FC8;
	tbl[878] = 15'h4FDB;
	tbl[879] = 15'h4FEF;
	tbl[880] = 15'h5003;
	tbl[881] = 15'h5016;
	tbl[882] = 15'h502A;
	tbl[883] = 15'h503E;
	tbl[884] = 15'h5051;
	tbl[885] = 15'h5065;
	tbl[886] = 15'h5078;
	tbl[887] = 15'h508C;
	tbl[888] = 15'h509F;
	tbl[889] = 15'h50B3;
	tbl[890] = 15'h50C6;
	tbl[891] = 15'h50DA;
	tbl[892] = 15'h50ED;
	tbl[893] = 15'h5101;
	tbl[894] = 15'h5114;
	tbl[895] = 15'h5128;
	tbl[896] = 15'h513B;
	tbl[897] = 15'h514F;
	tbl[898] = 15'h5162;
	tbl[899] = 15'h5175;
	tbl[900] = 15'h5189;
	tbl[901] = 15'h519C;
	tbl[902] = 15'h51B0;
	tbl[903] = 15'h51C3;
	tbl[904] = 15'h51D6;
	tbl[905] = 15'h51EA;
	tbl[906] = 15'h51FD;
	tbl[907] = 15'h5210;
	tbl[908] = 15'h5223;
	tbl[909] = 15'h5237;
	tbl[910] = 15'h524A;
	tbl[911] = 15'h525D;
	tbl[912] = 15'h5270;
	tbl[913] = 15'h5284;
	tbl[914] = 15'h5297;
	tbl[915] = 15'h52AA;
	tbl[916] = 15'h52BD;
	tbl[917] = 15'h52D1;
	tbl[918] = 15'h52E4;
	tbl[919] = 15'h52F7;
	tbl[920] = 15'h530A;
	tbl[921] = 15'h531D;
	tbl[922] = 15'h5330;
	tbl[923] = 15'h5343;
	tbl[924] = 15'h5356;
	tbl[925] = 15'h5369;
	tbl[926] = 15'h537D;
	tbl[927] = 15'h5390;
	tbl[928] = 15'h53A3;
	tbl[929] = 15'h53B6;
	tbl[930] = 15'h53C9;
	tbl[931] = 15'h53DC;
	tbl[932] = 15'h53EF;
	tbl[933] = 15'h5402;
	tbl[934] = 15'h5415;
	tbl[935] = 15'h5428;
	tbl[936] = 15'h543B;
	tbl[937] = 15'h544D;
	tbl[938] = 15'h5460;
	tbl[939] = 15'h5473;
	tbl[940] = 15'h5486;
	tbl[941] = 15'h5499;
	tbl[942] = 15'h54AC;
	tbl[943] = 15'h54BF;
	tbl[944] = 15'h54D2;
	tbl[945] = 15'h54E4;
	tbl[946] = 15'h54F7;
	tbl[947] = 15'h550A;
	tbl[948] = 15'h551D;
	tbl[949] = 15'h5530;
	tbl[950] = 15'h5542;
	tbl[951] = 15'h5555;
	tbl[952] = 15'h5568;
	tbl[953] = 15'h557B;
	tbl[954] = 15'h558D;
	tbl[955] = 15'h55A0;
	tbl[956] = 15'h55B3;
	tbl[957] = 15'h55C5;
	tbl[958] = 15'h55D8;
	tbl[959] = 15'h55EB;
	tbl[960] = 15'h55FD;
	tbl[961] = 15'h5610;
	tbl[962] = 15'h5622;
	tbl[963] = 15'h5635;
	tbl[964] = 15'h5648;
	tbl[965] = 15'h565A;
	tbl[966] = 15'h566D;
	tbl[967] = 15'h567F;
	tbl[968] = 15'h5692;
	tbl[969] = 15'h56A4;
	tbl[970] = 15'h56B7;
	tbl[971] = 15'h56C9;
	tbl[972] = 15'h56DC;
	tbl[973] = 15'h56EE;
	tbl[974] = 15'h5701;
	tbl[975] = 15'h5713;
	tbl[976] = 15'h5726;
	tbl[977] = 15'h5738;
	tbl[978] = 15'h574A;
	tbl[979] = 15'h575D;
	tbl[980] = 15'h576F;
	tbl[981] = 15'h5781;
	tbl[982] = 15'h5794;
	tbl[983] = 15'h57A6;
	tbl[984] = 15'h57B8;
	tbl[985] = 15'h57CB;
	tbl[986] = 15'h57DD;
	tbl[987] = 15'h57EF;
	tbl[988] = 15'h5802;
	tbl[989] = 15'h5814;
	tbl[990] = 15'h5826;
	tbl[991] = 15'h5838;
	tbl[992] = 15'h584A;
	tbl[993] = 15'h585D;
	tbl[994] = 15'h586F;
	tbl[995] = 15'h5881;
	tbl[996] = 15'h5893;
	tbl[997] = 15'h58A5;
	tbl[998] = 15'h58B7;
	tbl[999] = 15'h58CA;
	tbl[1000] = 15'h58DC;
	tbl[1001] = 15'h58EE;
	tbl[1002] = 15'h5900;
	tbl[1003] = 15'h5912;
	tbl[1004] = 15'h5924;
	tbl[1005] = 15'h5936;
	tbl[1006] = 15'h5948;
	tbl[1007] = 15'h595A;
	tbl[1008] = 15'h596C;
	tbl[1009] = 15'h597E;
	tbl[1010] = 15'h5990;
	tbl[1011] = 15'h59A2;
	tbl[1012] = 15'h59B4;
	tbl[1013] = 15'h59C6;
	tbl[1014] = 15'h59D8;
	tbl[1015] = 15'h59EA;
	tbl[1016] = 15'h59FC;
	tbl[1017] = 15'h5A0D;
	tbl[1018] = 15'h5A1F;
	tbl[1019] = 15'h5A31;
	tbl[1020] = 15'h5A43;
	tbl[1021] = 15'h5A55;
	tbl[1022] = 15'h5A67;
	tbl[1023] = 15'h5A78;
	tbl[1024] = 15'h5A8A;
	tbl[1025] = 15'h5A9C;
	tbl[1026] = 15'h5AAE;
	tbl[1027] = 15'h5ABF;
	tbl[1028] = 15'h5AD1;
	tbl[1029] = 15'h5AE3;
	tbl[1030] = 15'h5AF5;
	tbl[1031] = 15'h5B06;
	tbl[1032] = 15'h5B18;
	tbl[1033] = 15'h5B2A;
	tbl[1034] = 15'h5B3B;
	tbl[1035] = 15'h5B4D;
	tbl[1036] = 15'h5B5E;
	tbl[1037] = 15'h5B70;
	tbl[1038] = 15'h5B82;
	tbl[1039] = 15'h5B93;
	tbl[1040] = 15'h5BA5;
	tbl[1041] = 15'h5BB6;
	tbl[1042] = 15'h5BC8;
	tbl[1043] = 15'h5BD9;
	tbl[1044] = 15'h5BEB;
	tbl[1045] = 15'h5BFC;
	tbl[1046] = 15'h5C0E;
	tbl[1047] = 15'h5C1F;
	tbl[1048] = 15'h5C31;
	tbl[1049] = 15'h5C42;
	tbl[1050] = 15'h5C54;
	tbl[1051] = 15'h5C65;
	tbl[1052] = 15'h5C76;
	tbl[1053] = 15'h5C88;
	tbl[1054] = 15'h5C99;
	tbl[1055] = 15'h5CAB;
	tbl[1056] = 15'h5CBC;
	tbl[1057] = 15'h5CCD;
	tbl[1058] = 15'h5CDE;
	tbl[1059] = 15'h5CF0;
	tbl[1060] = 15'h5D01;
	tbl[1061] = 15'h5D12;
	tbl[1062] = 15'h5D24;
	tbl[1063] = 15'h5D35;
	tbl[1064] = 15'h5D46;
	tbl[1065] = 15'h5D57;
	tbl[1066] = 15'h5D68;
	tbl[1067] = 15'h5D7A;
	tbl[1068] = 15'h5D8B;
	tbl[1069] = 15'h5D9C;
	tbl[1070] = 15'h5DAD;
	tbl[1071] = 15'h5DBE;
	tbl[1072] = 15'h5DCF;
	tbl[1073] = 15'h5DE0;
	tbl[1074] = 15'h5DF2;
	tbl[1075] = 15'h5E03;
	tbl[1076] = 15'h5E14;
	tbl[1077] = 15'h5E25;
	tbl[1078] = 15'h5E36;
	tbl[1079] = 15'h5E47;
	tbl[1080] = 15'h5E58;
	tbl[1081] = 15'h5E69;
	tbl[1082] = 15'h5E7A;
	tbl[1083] = 15'h5E8B;
	tbl[1084] = 15'h5E9C;
	tbl[1085] = 15'h5EAD;
	tbl[1086] = 15'h5EBD;
	tbl[1087] = 15'h5ECE;
	tbl[1088] = 15'h5EDF;
	tbl[1089] = 15'h5EF0;
	tbl[1090] = 15'h5F01;
	tbl[1091] = 15'h5F12;
	tbl[1092] = 15'h5F23;
	tbl[1093] = 15'h5F33;
	tbl[1094] = 15'h5F44;
	tbl[1095] = 15'h5F55;
	tbl[1096] = 15'h5F66;
	tbl[1097] = 15'h5F77;
	tbl[1098] = 15'h5F87;
	tbl[1099] = 15'h5F98;
	tbl[1100] = 15'h5FA9;
	tbl[1101] = 15'h5FB9;
	tbl[1102] = 15'h5FCA;
	tbl[1103] = 15'h5FDB;
	tbl[1104] = 15'h5FEB;
	tbl[1105] = 15'h5FFC;
	tbl[1106] = 15'h600D;
	tbl[1107] = 15'h601D;
	tbl[1108] = 15'h602E;
	tbl[1109] = 15'h603E;
	tbl[1110] = 15'h604F;
	tbl[1111] = 15'h6060;
	tbl[1112] = 15'h6070;
	tbl[1113] = 15'h6081;
	tbl[1114] = 15'h6091;
	tbl[1115] = 15'h60A2;
	tbl[1116] = 15'h60B2;
	tbl[1117] = 15'h60C3;
	tbl[1118] = 15'h60D3;
	tbl[1119] = 15'h60E4;
	tbl[1120] = 15'h60F4;
	tbl[1121] = 15'h6104;
	tbl[1122] = 15'h6115;
	tbl[1123] = 15'h6125;
	tbl[1124] = 15'h6135;
	tbl[1125] = 15'h6146;
	tbl[1126] = 15'h6156;
	tbl[1127] = 15'h6166;
	tbl[1128] = 15'h6177;
	tbl[1129] = 15'h6187;
	tbl[1130] = 15'h6197;
	tbl[1131] = 15'h61A8;
	tbl[1132] = 15'h61B8;
	tbl[1133] = 15'h61C8;
	tbl[1134] = 15'h61D8;
	tbl[1135] = 15'h61E9;
	tbl[1136] = 15'h61F9;
	tbl[1137] = 15'h6209;
	tbl[1138] = 15'h6219;
	tbl[1139] = 15'h6229;
	tbl[1140] = 15'h6239;
	tbl[1141] = 15'h6249;
	tbl[1142] = 15'h625A;
	tbl[1143] = 15'h626A;
	tbl[1144] = 15'h627A;
	tbl[1145] = 15'h628A;
	tbl[1146] = 15'h629A;
	tbl[1147] = 15'h62AA;
	tbl[1148] = 15'h62BA;
	tbl[1149] = 15'h62CA;
	tbl[1150] = 15'h62DA;
	tbl[1151] = 15'h62EA;
	tbl[1152] = 15'h62FA;
	tbl[1153] = 15'h630A;
	tbl[1154] = 15'h631A;
	tbl[1155] = 15'h6329;
	tbl[1156] = 15'h6339;
	tbl[1157] = 15'h6349;
	tbl[1158] = 15'h6359;
	tbl[1159] = 15'h6369;
	tbl[1160] = 15'h6379;
	tbl[1161] = 15'h6389;
	tbl[1162] = 15'h6398;
	tbl[1163] = 15'h63A8;
	tbl[1164] = 15'h63B8;
	tbl[1165] = 15'h63C8;
	tbl[1166] = 15'h63D7;
	tbl[1167] = 15'h63E7;
	tbl[1168] = 15'h63F7;
	tbl[1169] = 15'h6407;
	tbl[1170] = 15'h6416;
	tbl[1171] = 15'h6426;
	tbl[1172] = 15'h6436;
	tbl[1173] = 15'h6445;
	tbl[1174] = 15'h6455;
	tbl[1175] = 15'h6464;
	tbl[1176] = 15'h6474;
	tbl[1177] = 15'h6484;
	tbl[1178] = 15'h6493;
	tbl[1179] = 15'h64A3;
	tbl[1180] = 15'h64B2;
	tbl[1181] = 15'h64C2;
	tbl[1182] = 15'h64D1;
	tbl[1183] = 15'h64E1;
	tbl[1184] = 15'h64F0;
	tbl[1185] = 15'h6500;
	tbl[1186] = 15'h650F;
	tbl[1187] = 15'h651F;
	tbl[1188] = 15'h652E;
	tbl[1189] = 15'h653D;
	tbl[1190] = 15'h654D;
	tbl[1191] = 15'h655C;
	tbl[1192] = 15'h656B;
	tbl[1193] = 15'h657B;
	tbl[1194] = 15'h658A;
	tbl[1195] = 15'h6599;
	tbl[1196] = 15'h65A9;
	tbl[1197] = 15'h65B8;
	tbl[1198] = 15'h65C7;
	tbl[1199] = 15'h65D6;
	tbl[1200] = 15'h65E6;
	tbl[1201] = 15'h65F5;
	tbl[1202] = 15'h6604;
	tbl[1203] = 15'h6613;
	tbl[1204] = 15'h6622;
	tbl[1205] = 15'h6631;
	tbl[1206] = 15'h6641;
	tbl[1207] = 15'h6650;
	tbl[1208] = 15'h665F;
	tbl[1209] = 15'h666E;
	tbl[1210] = 15'h667D;
	tbl[1211] = 15'h668C;
	tbl[1212] = 15'h669B;
	tbl[1213] = 15'h66AA;
	tbl[1214] = 15'h66B9;
	tbl[1215] = 15'h66C8;
	tbl[1216] = 15'h66D7;
	tbl[1217] = 15'h66E6;
	tbl[1218] = 15'h66F5;
	tbl[1219] = 15'h6704;
	tbl[1220] = 15'h6713;
	tbl[1221] = 15'h6722;
	tbl[1222] = 15'h6731;
	tbl[1223] = 15'h673F;
	tbl[1224] = 15'h674E;
	tbl[1225] = 15'h675D;
	tbl[1226] = 15'h676C;
	tbl[1227] = 15'h677B;
	tbl[1228] = 15'h678A;
	tbl[1229] = 15'h6798;
	tbl[1230] = 15'h67A7;
	tbl[1231] = 15'h67B6;
	tbl[1232] = 15'h67C5;
	tbl[1233] = 15'h67D3;
	tbl[1234] = 15'h67E2;
	tbl[1235] = 15'h67F1;
	tbl[1236] = 15'h67FF;
	tbl[1237] = 15'h680E;
	tbl[1238] = 15'h681D;
	tbl[1239] = 15'h682B;
	tbl[1240] = 15'h683A;
	tbl[1241] = 15'h6848;
	tbl[1242] = 15'h6857;
	tbl[1243] = 15'h6866;
	tbl[1244] = 15'h6874;
	tbl[1245] = 15'h6883;
	tbl[1246] = 15'h6891;
	tbl[1247] = 15'h68A0;
	tbl[1248] = 15'h68AE;
	tbl[1249] = 15'h68BD;
	tbl[1250] = 15'h68CB;
	tbl[1251] = 15'h68D9;
	tbl[1252] = 15'h68E8;
	tbl[1253] = 15'h68F6;
	tbl[1254] = 15'h6905;
	tbl[1255] = 15'h6913;
	tbl[1256] = 15'h6921;
	tbl[1257] = 15'h6930;
	tbl[1258] = 15'h693E;
	tbl[1259] = 15'h694C;
	tbl[1260] = 15'h695B;
	tbl[1261] = 15'h6969;
	tbl[1262] = 15'h6977;
	tbl[1263] = 15'h6985;
	tbl[1264] = 15'h6994;
	tbl[1265] = 15'h69A2;
	tbl[1266] = 15'h69B0;
	tbl[1267] = 15'h69BE;
	tbl[1268] = 15'h69CC;
	tbl[1269] = 15'h69DA;
	tbl[1270] = 15'h69E9;
	tbl[1271] = 15'h69F7;
	tbl[1272] = 15'h6A05;
	tbl[1273] = 15'h6A13;
	tbl[1274] = 15'h6A21;
	tbl[1275] = 15'h6A2F;
	tbl[1276] = 15'h6A3D;
	tbl[1277] = 15'h6A4B;
	tbl[1278] = 15'h6A59;
	tbl[1279] = 15'h6A67;
	tbl[1280] = 15'h6A75;
	tbl[1281] = 15'h6A83;
	tbl[1282] = 15'h6A91;
	tbl[1283] = 15'h6A9F;
	tbl[1284] = 15'h6AAD;
	tbl[1285] = 15'h6ABB;
	tbl[1286] = 15'h6AC8;
	tbl[1287] = 15'h6AD6;
	tbl[1288] = 15'h6AE4;
	tbl[1289] = 15'h6AF2;
	tbl[1290] = 15'h6B00;
	tbl[1291] = 15'h6B0E;
	tbl[1292] = 15'h6B1B;
	tbl[1293] = 15'h6B29;
	tbl[1294] = 15'h6B37;
	tbl[1295] = 15'h6B45;
	tbl[1296] = 15'h6B52;
	tbl[1297] = 15'h6B60;
	tbl[1298] = 15'h6B6E;
	tbl[1299] = 15'h6B7B;
	tbl[1300] = 15'h6B89;
	tbl[1301] = 15'h6B97;
	tbl[1302] = 15'h6BA4;
	tbl[1303] = 15'h6BB2;
	tbl[1304] = 15'h6BBF;
	tbl[1305] = 15'h6BCD;
	tbl[1306] = 15'h6BDA;
	tbl[1307] = 15'h6BE8;
	tbl[1308] = 15'h6BF6;
	tbl[1309] = 15'h6C03;
	tbl[1310] = 15'h6C11;
	tbl[1311] = 15'h6C1E;
	tbl[1312] = 15'h6C2B;
	tbl[1313] = 15'h6C39;
	tbl[1314] = 15'h6C46;
	tbl[1315] = 15'h6C54;
	tbl[1316] = 15'h6C61;
	tbl[1317] = 15'h6C6E;
	tbl[1318] = 15'h6C7C;
	tbl[1319] = 15'h6C89;
	tbl[1320] = 15'h6C96;
	tbl[1321] = 15'h6CA4;
	tbl[1322] = 15'h6CB1;
	tbl[1323] = 15'h6CBE;
	tbl[1324] = 15'h6CCC;
	tbl[1325] = 15'h6CD9;
	tbl[1326] = 15'h6CE6;
	tbl[1327] = 15'h6CF3;
	tbl[1328] = 15'h6D00;
	tbl[1329] = 15'h6D0E;
	tbl[1330] = 15'h6D1B;
	tbl[1331] = 15'h6D28;
	tbl[1332] = 15'h6D35;
	tbl[1333] = 15'h6D42;
	tbl[1334] = 15'h6D4F;
	tbl[1335] = 15'h6D5C;
	tbl[1336] = 15'h6D69;
	tbl[1337] = 15'h6D76;
	tbl[1338] = 15'h6D83;
	tbl[1339] = 15'h6D90;
	tbl[1340] = 15'h6D9D;
	tbl[1341] = 15'h6DAA;
	tbl[1342] = 15'h6DB7;
	tbl[1343] = 15'h6DC4;
	tbl[1344] = 15'h6DD1;
	tbl[1345] = 15'h6DDE;
	tbl[1346] = 15'h6DEB;
	tbl[1347] = 15'h6DF8;
	tbl[1348] = 15'h6E05;
	tbl[1349] = 15'h6E12;
	tbl[1350] = 15'h6E1E;
	tbl[1351] = 15'h6E2B;
	tbl[1352] = 15'h6E38;
	tbl[1353] = 15'h6E45;
	tbl[1354] = 15'h6E52;
	tbl[1355] = 15'h6E5E;
	tbl[1356] = 15'h6E6B;
	tbl[1357] = 15'h6E78;
	tbl[1358] = 15'h6E84;
	tbl[1359] = 15'h6E91;
	tbl[1360] = 15'h6E9E;
	tbl[1361] = 15'h6EAA;
	tbl[1362] = 15'h6EB7;
	tbl[1363] = 15'h6EC4;
	tbl[1364] = 15'h6ED0;
	tbl[1365] = 15'h6EDD;
	tbl[1366] = 15'h6EE9;
	tbl[1367] = 15'h6EF6;
	tbl[1368] = 15'h6F02;
	tbl[1369] = 15'h6F0F;
	tbl[1370] = 15'h6F1B;
	tbl[1371] = 15'h6F28;
	tbl[1372] = 15'h6F34;
	tbl[1373] = 15'h6F41;
	tbl[1374] = 15'h6F4D;
	tbl[1375] = 15'h6F5A;
	tbl[1376] = 15'h6F66;
	tbl[1377] = 15'h6F72;
	tbl[1378] = 15'h6F7F;
	tbl[1379] = 15'h6F8B;
	tbl[1380] = 15'h6F97;
	tbl[1381] = 15'h6FA4;
	tbl[1382] = 15'h6FB0;
	tbl[1383] = 15'h6FBC;
	tbl[1384] = 15'h6FC8;
	tbl[1385] = 15'h6FD5;
	tbl[1386] = 15'h6FE1;
	tbl[1387] = 15'h6FED;
	tbl[1388] = 15'h6FF9;
	tbl[1389] = 15'h7006;
	tbl[1390] = 15'h7012;
	tbl[1391] = 15'h701E;
	tbl[1392] = 15'h702A;
	tbl[1393] = 15'h7036;
	tbl[1394] = 15'h7042;
	tbl[1395] = 15'h704E;
	tbl[1396] = 15'h705A;
	tbl[1397] = 15'h7066;
	tbl[1398] = 15'h7072;
	tbl[1399] = 15'h707E;
	tbl[1400] = 15'h708A;
	tbl[1401] = 15'h7096;
	tbl[1402] = 15'h70A2;
	tbl[1403] = 15'h70AE;
	tbl[1404] = 15'h70BA;
	tbl[1405] = 15'h70C6;
	tbl[1406] = 15'h70D2;
	tbl[1407] = 15'h70DE;
	tbl[1408] = 15'h70EA;
	tbl[1409] = 15'h70F5;
	tbl[1410] = 15'h7101;
	tbl[1411] = 15'h710D;
	tbl[1412] = 15'h7119;
	tbl[1413] = 15'h7125;
	tbl[1414] = 15'h7130;
	tbl[1415] = 15'h713C;
	tbl[1416] = 15'h7148;
	tbl[1417] = 15'h7153;
	tbl[1418] = 15'h715F;
	tbl[1419] = 15'h716B;
	tbl[1420] = 15'h7176;
	tbl[1421] = 15'h7182;
	tbl[1422] = 15'h718E;
	tbl[1423] = 15'h7199;
	tbl[1424] = 15'h71A5;
	tbl[1425] = 15'h71B0;
	tbl[1426] = 15'h71BC;
	tbl[1427] = 15'h71C7;
	tbl[1428] = 15'h71D3;
	tbl[1429] = 15'h71DE;
	tbl[1430] = 15'h71EA;
	tbl[1431] = 15'h71F5;
	tbl[1432] = 15'h7201;
	tbl[1433] = 15'h720C;
	tbl[1434] = 15'h7218;
	tbl[1435] = 15'h7223;
	tbl[1436] = 15'h722E;
	tbl[1437] = 15'h723A;
	tbl[1438] = 15'h7245;
	tbl[1439] = 15'h7250;
	tbl[1440] = 15'h725C;
	tbl[1441] = 15'h7267;
	tbl[1442] = 15'h7272;
	tbl[1443] = 15'h727E;
	tbl[1444] = 15'h7289;
	tbl[1445] = 15'h7294;
	tbl[1446] = 15'h729F;
	tbl[1447] = 15'h72AA;
	tbl[1448] = 15'h72B6;
	tbl[1449] = 15'h72C1;
	tbl[1450] = 15'h72CC;
	tbl[1451] = 15'h72D7;
	tbl[1452] = 15'h72E2;
	tbl[1453] = 15'h72ED;
	tbl[1454] = 15'h72F8;
	tbl[1455] = 15'h7303;
	tbl[1456] = 15'h730E;
	tbl[1457] = 15'h7319;
	tbl[1458] = 15'h7324;
	tbl[1459] = 15'h732F;
	tbl[1460] = 15'h733A;
	tbl[1461] = 15'h7345;
	tbl[1462] = 15'h7350;
	tbl[1463] = 15'h735B;
	tbl[1464] = 15'h7366;
	tbl[1465] = 15'h7371;
	tbl[1466] = 15'h737B;
	tbl[1467] = 15'h7386;
	tbl[1468] = 15'h7391;
	tbl[1469] = 15'h739C;
	tbl[1470] = 15'h73A7;
	tbl[1471] = 15'h73B1;
	tbl[1472] = 15'h73BC;
	tbl[1473] = 15'h73C7;
	tbl[1474] = 15'h73D2;
	tbl[1475] = 15'h73DC;
	tbl[1476] = 15'h73E7;
	tbl[1477] = 15'h73F2;
	tbl[1478] = 15'h73FC;
	tbl[1479] = 15'h7407;
	tbl[1480] = 15'h7412;
	tbl[1481] = 15'h741C;
	tbl[1482] = 15'h7427;
	tbl[1483] = 15'h7431;
	tbl[1484] = 15'h743C;
	tbl[1485] = 15'h7446;
	tbl[1486] = 15'h7451;
	tbl[1487] = 15'h745B;
	tbl[1488] = 15'h7466;
	tbl[1489] = 15'h7470;
	tbl[1490] = 15'h747B;
	tbl[1491] = 15'h7485;
	tbl[1492] = 15'h7490;
	tbl[1493] = 15'h749A;
	tbl[1494] = 15'h74A4;
	tbl[1495] = 15'h74AF;
	tbl[1496] = 15'h74B9;
	tbl[1497] = 15'h74C3;
	tbl[1498] = 15'h74CE;
	tbl[1499] = 15'h74D8;
	tbl[1500] = 15'h74E2;
	tbl[1501] = 15'h74EC;
	tbl[1502] = 15'h74F7;
	tbl[1503] = 15'h7501;
	tbl[1504] = 15'h750B;
	tbl[1505] = 15'h7515;
	tbl[1506] = 15'h751F;
	tbl[1507] = 15'h7529;
	tbl[1508] = 15'h7533;
	tbl[1509] = 15'h753E;
	tbl[1510] = 15'h7548;
	tbl[1511] = 15'h7552;
	tbl[1512] = 15'h755C;
	tbl[1513] = 15'h7566;
	tbl[1514] = 15'h7570;
	tbl[1515] = 15'h757A;
	tbl[1516] = 15'h7584;
	tbl[1517] = 15'h758E;
	tbl[1518] = 15'h7598;
	tbl[1519] = 15'h75A2;
	tbl[1520] = 15'h75AB;
	tbl[1521] = 15'h75B5;
	tbl[1522] = 15'h75BF;
	tbl[1523] = 15'h75C9;
	tbl[1524] = 15'h75D3;
	tbl[1525] = 15'h75DD;
	tbl[1526] = 15'h75E6;
	tbl[1527] = 15'h75F0;
	tbl[1528] = 15'h75FA;
	tbl[1529] = 15'h7604;
	tbl[1530] = 15'h760D;
	tbl[1531] = 15'h7617;
	tbl[1532] = 15'h7621;
	tbl[1533] = 15'h762B;
	tbl[1534] = 15'h7634;
	tbl[1535] = 15'h763E;
	tbl[1536] = 15'h7647;
	tbl[1537] = 15'h7651;
	tbl[1538] = 15'h765B;
	tbl[1539] = 15'h7664;
	tbl[1540] = 15'h766E;
	tbl[1541] = 15'h7677;
	tbl[1542] = 15'h7681;
	tbl[1543] = 15'h768A;
	tbl[1544] = 15'h7694;
	tbl[1545] = 15'h769D;
	tbl[1546] = 15'h76A7;
	tbl[1547] = 15'h76B0;
	tbl[1548] = 15'h76B9;
	tbl[1549] = 15'h76C3;
	tbl[1550] = 15'h76CC;
	tbl[1551] = 15'h76D6;
	tbl[1552] = 15'h76DF;
	tbl[1553] = 15'h76E8;
	tbl[1554] = 15'h76F2;
	tbl[1555] = 15'h76FB;
	tbl[1556] = 15'h7704;
	tbl[1557] = 15'h770D;
	tbl[1558] = 15'h7717;
	tbl[1559] = 15'h7720;
	tbl[1560] = 15'h7729;
	tbl[1561] = 15'h7732;
	tbl[1562] = 15'h773B;
	tbl[1563] = 15'h7744;
	tbl[1564] = 15'h774E;
	tbl[1565] = 15'h7757;
	tbl[1566] = 15'h7760;
	tbl[1567] = 15'h7769;
	tbl[1568] = 15'h7772;
	tbl[1569] = 15'h777B;
	tbl[1570] = 15'h7784;
	tbl[1571] = 15'h778D;
	tbl[1572] = 15'h7796;
	tbl[1573] = 15'h779F;
	tbl[1574] = 15'h77A8;
	tbl[1575] = 15'h77B1;
	tbl[1576] = 15'h77BA;
	tbl[1577] = 15'h77C2;
	tbl[1578] = 15'h77CB;
	tbl[1579] = 15'h77D4;
	tbl[1580] = 15'h77DD;
	tbl[1581] = 15'h77E6;
	tbl[1582] = 15'h77EF;
	tbl[1583] = 15'h77F7;
	tbl[1584] = 15'h7800;
	tbl[1585] = 15'h7809;
	tbl[1586] = 15'h7812;
	tbl[1587] = 15'h781A;
	tbl[1588] = 15'h7823;
	tbl[1589] = 15'h782C;
	tbl[1590] = 15'h7834;
	tbl[1591] = 15'h783D;
	tbl[1592] = 15'h7845;
	tbl[1593] = 15'h784E;
	tbl[1594] = 15'h7857;
	tbl[1595] = 15'h785F;
	tbl[1596] = 15'h7868;
	tbl[1597] = 15'h7870;
	tbl[1598] = 15'h7879;
	tbl[1599] = 15'h7881;
	tbl[1600] = 15'h788A;
	tbl[1601] = 15'h7892;
	tbl[1602] = 15'h789B;
	tbl[1603] = 15'h78A3;
	tbl[1604] = 15'h78AB;
	tbl[1605] = 15'h78B4;
	tbl[1606] = 15'h78BC;
	tbl[1607] = 15'h78C4;
	tbl[1608] = 15'h78CD;
	tbl[1609] = 15'h78D5;
	tbl[1610] = 15'h78DD;
	tbl[1611] = 15'h78E6;
	tbl[1612] = 15'h78EE;
	tbl[1613] = 15'h78F6;
	tbl[1614] = 15'h78FE;
	tbl[1615] = 15'h7906;
	tbl[1616] = 15'h790F;
	tbl[1617] = 15'h7917;
	tbl[1618] = 15'h791F;
	tbl[1619] = 15'h7927;
	tbl[1620] = 15'h792F;
	tbl[1621] = 15'h7937;
	tbl[1622] = 15'h793F;
	tbl[1623] = 15'h7947;
	tbl[1624] = 15'h794F;
	tbl[1625] = 15'h7957;
	tbl[1626] = 15'h795F;
	tbl[1627] = 15'h7967;
	tbl[1628] = 15'h796F;
	tbl[1629] = 15'h7977;
	tbl[1630] = 15'h797F;
	tbl[1631] = 15'h7987;
	tbl[1632] = 15'h798F;
	tbl[1633] = 15'h7997;
	tbl[1634] = 15'h799F;
	tbl[1635] = 15'h79A7;
	tbl[1636] = 15'h79AE;
	tbl[1637] = 15'h79B6;
	tbl[1638] = 15'h79BE;
	tbl[1639] = 15'h79C6;
	tbl[1640] = 15'h79CD;
	tbl[1641] = 15'h79D5;
	tbl[1642] = 15'h79DD;
	tbl[1643] = 15'h79E4;
	tbl[1644] = 15'h79EC;
	tbl[1645] = 15'h79F4;
	tbl[1646] = 15'h79FB;
	tbl[1647] = 15'h7A03;
	tbl[1648] = 15'h7A0B;
	tbl[1649] = 15'h7A12;
	tbl[1650] = 15'h7A1A;
	tbl[1651] = 15'h7A21;
	tbl[1652] = 15'h7A29;
	tbl[1653] = 15'h7A30;
	tbl[1654] = 15'h7A38;
	tbl[1655] = 15'h7A3F;
	tbl[1656] = 15'h7A47;
	tbl[1657] = 15'h7A4E;
	tbl[1658] = 15'h7A55;
	tbl[1659] = 15'h7A5D;
	tbl[1660] = 15'h7A64;
	tbl[1661] = 15'h7A6C;
	tbl[1662] = 15'h7A73;
	tbl[1663] = 15'h7A7A;
	tbl[1664] = 15'h7A81;
	tbl[1665] = 15'h7A89;
	tbl[1666] = 15'h7A90;
	tbl[1667] = 15'h7A97;
	tbl[1668] = 15'h7A9E;
	tbl[1669] = 15'h7AA6;
	tbl[1670] = 15'h7AAD;
	tbl[1671] = 15'h7AB4;
	tbl[1672] = 15'h7ABB;
	tbl[1673] = 15'h7AC2;
	tbl[1674] = 15'h7AC9;
	tbl[1675] = 15'h7AD0;
	tbl[1676] = 15'h7AD8;
	tbl[1677] = 15'h7ADF;
	tbl[1678] = 15'h7AE6;
	tbl[1679] = 15'h7AED;
	tbl[1680] = 15'h7AF4;
	tbl[1681] = 15'h7AFB;
	tbl[1682] = 15'h7B02;
	tbl[1683] = 15'h7B09;
	tbl[1684] = 15'h7B0F;
	tbl[1685] = 15'h7B16;
	tbl[1686] = 15'h7B1D;
	tbl[1687] = 15'h7B24;
	tbl[1688] = 15'h7B2B;
	tbl[1689] = 15'h7B32;
	tbl[1690] = 15'h7B39;
	tbl[1691] = 15'h7B3F;
	tbl[1692] = 15'h7B46;
	tbl[1693] = 15'h7B4D;
	tbl[1694] = 15'h7B54;
	tbl[1695] = 15'h7B5A;
	tbl[1696] = 15'h7B61;
	tbl[1697] = 15'h7B68;
	tbl[1698] = 15'h7B6E;
	tbl[1699] = 15'h7B75;
	tbl[1700] = 15'h7B7C;
	tbl[1701] = 15'h7B82;
	tbl[1702] = 15'h7B89;
	tbl[1703] = 15'h7B8F;
	tbl[1704] = 15'h7B96;
	tbl[1705] = 15'h7B9D;
	tbl[1706] = 15'h7BA3;
	tbl[1707] = 15'h7BAA;
	tbl[1708] = 15'h7BB0;
	tbl[1709] = 15'h7BB7;
	tbl[1710] = 15'h7BBD;
	tbl[1711] = 15'h7BC3;
	tbl[1712] = 15'h7BCA;
	tbl[1713] = 15'h7BD0;
	tbl[1714] = 15'h7BD7;
	tbl[1715] = 15'h7BDD;
	tbl[1716] = 15'h7BE3;
	tbl[1717] = 15'h7BE9;
	tbl[1718] = 15'h7BF0;
	tbl[1719] = 15'h7BF6;
	tbl[1720] = 15'h7BFC;
	tbl[1721] = 15'h7C03;
	tbl[1722] = 15'h7C09;
	tbl[1723] = 15'h7C0F;
	tbl[1724] = 15'h7C15;
	tbl[1725] = 15'h7C1B;
	tbl[1726] = 15'h7C21;
	tbl[1727] = 15'h7C28;
	tbl[1728] = 15'h7C2E;
	tbl[1729] = 15'h7C34;
	tbl[1730] = 15'h7C3A;
	tbl[1731] = 15'h7C40;
	tbl[1732] = 15'h7C46;
	tbl[1733] = 15'h7C4C;
	tbl[1734] = 15'h7C52;
	tbl[1735] = 15'h7C58;
	tbl[1736] = 15'h7C5E;
	tbl[1737] = 15'h7C64;
	tbl[1738] = 15'h7C6A;
	tbl[1739] = 15'h7C70;
	tbl[1740] = 15'h7C75;
	tbl[1741] = 15'h7C7B;
	tbl[1742] = 15'h7C81;
	tbl[1743] = 15'h7C87;
	tbl[1744] = 15'h7C8D;
	tbl[1745] = 15'h7C93;
	tbl[1746] = 15'h7C98;
	tbl[1747] = 15'h7C9E;
	tbl[1748] = 15'h7CA4;
	tbl[1749] = 15'h7CA9;
	tbl[1750] = 15'h7CAF;
	tbl[1751] = 15'h7CB5;
	tbl[1752] = 15'h7CBB;
	tbl[1753] = 15'h7CC0;
	tbl[1754] = 15'h7CC6;
	tbl[1755] = 15'h7CCB;
	tbl[1756] = 15'h7CD1;
	tbl[1757] = 15'h7CD6;
	tbl[1758] = 15'h7CDC;
	tbl[1759] = 15'h7CE2;
	tbl[1760] = 15'h7CE7;
	tbl[1761] = 15'h7CED;
	tbl[1762] = 15'h7CF2;
	tbl[1763] = 15'h7CF7;
	tbl[1764] = 15'h7CFD;
	tbl[1765] = 15'h7D02;
	tbl[1766] = 15'h7D08;
	tbl[1767] = 15'h7D0D;
	tbl[1768] = 15'h7D12;
	tbl[1769] = 15'h7D18;
	tbl[1770] = 15'h7D1D;
	tbl[1771] = 15'h7D22;
	tbl[1772] = 15'h7D28;
	tbl[1773] = 15'h7D2D;
	tbl[1774] = 15'h7D32;
	tbl[1775] = 15'h7D37;
	tbl[1776] = 15'h7D3D;
	tbl[1777] = 15'h7D42;
	tbl[1778] = 15'h7D47;
	tbl[1779] = 15'h7D4C;
	tbl[1780] = 15'h7D51;
	tbl[1781] = 15'h7D56;
	tbl[1782] = 15'h7D5B;
	tbl[1783] = 15'h7D60;
	tbl[1784] = 15'h7D65;
	tbl[1785] = 15'h7D6A;
	tbl[1786] = 15'h7D70;
	tbl[1787] = 15'h7D74;
	tbl[1788] = 15'h7D79;
	tbl[1789] = 15'h7D7E;
	tbl[1790] = 15'h7D83;
	tbl[1791] = 15'h7D88;
	tbl[1792] = 15'h7D8D;
	tbl[1793] = 15'h7D92;
	tbl[1794] = 15'h7D97;
	tbl[1795] = 15'h7D9C;
	tbl[1796] = 15'h7DA1;
	tbl[1797] = 15'h7DA5;
	tbl[1798] = 15'h7DAA;
	tbl[1799] = 15'h7DAF;
	tbl[1800] = 15'h7DB4;
	tbl[1801] = 15'h7DB8;
	tbl[1802] = 15'h7DBD;
	tbl[1803] = 15'h7DC2;
	tbl[1804] = 15'h7DC6;
	tbl[1805] = 15'h7DCB;
	tbl[1806] = 15'h7DD0;
	tbl[1807] = 15'h7DD4;
	tbl[1808] = 15'h7DD9;
	tbl[1809] = 15'h7DDE;
	tbl[1810] = 15'h7DE2;
	tbl[1811] = 15'h7DE7;
	tbl[1812] = 15'h7DEB;
	tbl[1813] = 15'h7DF0;
	tbl[1814] = 15'h7DF4;
	tbl[1815] = 15'h7DF9;
	tbl[1816] = 15'h7DFD;
	tbl[1817] = 15'h7E01;
	tbl[1818] = 15'h7E06;
	tbl[1819] = 15'h7E0A;
	tbl[1820] = 15'h7E0F;
	tbl[1821] = 15'h7E13;
	tbl[1822] = 15'h7E17;
	tbl[1823] = 15'h7E1C;
	tbl[1824] = 15'h7E20;
	tbl[1825] = 15'h7E24;
	tbl[1826] = 15'h7E28;
	tbl[1827] = 15'h7E2D;
	tbl[1828] = 15'h7E31;
	tbl[1829] = 15'h7E35;
	tbl[1830] = 15'h7E39;
	tbl[1831] = 15'h7E3D;
	tbl[1832] = 15'h7E42;
	tbl[1833] = 15'h7E46;
	tbl[1834] = 15'h7E4A;
	tbl[1835] = 15'h7E4E;
	tbl[1836] = 15'h7E52;
	tbl[1837] = 15'h7E56;
	tbl[1838] = 15'h7E5A;
	tbl[1839] = 15'h7E5E;
	tbl[1840] = 15'h7E62;
	tbl[1841] = 15'h7E66;
	tbl[1842] = 15'h7E6A;
	tbl[1843] = 15'h7E6E;
	tbl[1844] = 15'h7E72;
	tbl[1845] = 15'h7E76;
	tbl[1846] = 15'h7E7A;
	tbl[1847] = 15'h7E7D;
	tbl[1848] = 15'h7E81;
	tbl[1849] = 15'h7E85;
	tbl[1850] = 15'h7E89;
	tbl[1851] = 15'h7E8D;
	tbl[1852] = 15'h7E90;
	tbl[1853] = 15'h7E94;
	tbl[1854] = 15'h7E98;
	tbl[1855] = 15'h7E9C;
	tbl[1856] = 15'h7E9F;
	tbl[1857] = 15'h7EA3;
	tbl[1858] = 15'h7EA6;
	tbl[1859] = 15'h7EAA;
	tbl[1860] = 15'h7EAE;
	tbl[1861] = 15'h7EB1;
	tbl[1862] = 15'h7EB5;
	tbl[1863] = 15'h7EB8;
	tbl[1864] = 15'h7EBC;
	tbl[1865] = 15'h7EBF;
	tbl[1866] = 15'h7EC3;
	tbl[1867] = 15'h7EC6;
	tbl[1868] = 15'h7ECA;
	tbl[1869] = 15'h7ECD;
	tbl[1870] = 15'h7ED1;
	tbl[1871] = 15'h7ED4;
	tbl[1872] = 15'h7ED7;
	tbl[1873] = 15'h7EDB;
	tbl[1874] = 15'h7EDE;
	tbl[1875] = 15'h7EE2;
	tbl[1876] = 15'h7EE5;
	tbl[1877] = 15'h7EE8;
	tbl[1878] = 15'h7EEB;
	tbl[1879] = 15'h7EEF;
	tbl[1880] = 15'h7EF2;
	tbl[1881] = 15'h7EF5;
	tbl[1882] = 15'h7EF8;
	tbl[1883] = 15'h7EFB;
	tbl[1884] = 15'h7EFF;
	tbl[1885] = 15'h7F02;
	tbl[1886] = 15'h7F05;
	tbl[1887] = 15'h7F08;
	tbl[1888] = 15'h7F0B;
	tbl[1889] = 15'h7F0E;
	tbl[1890] = 15'h7F11;
	tbl[1891] = 15'h7F14;
	tbl[1892] = 15'h7F17;
	tbl[1893] = 15'h7F1A;
	tbl[1894] = 15'h7F1D;
	tbl[1895] = 15'h7F20;
	tbl[1896] = 15'h7F23;
	tbl[1897] = 15'h7F26;
	tbl[1898] = 15'h7F29;
	tbl[1899] = 15'h7F2B;
	tbl[1900] = 15'h7F2E;
	tbl[1901] = 15'h7F31;
	tbl[1902] = 15'h7F34;
	tbl[1903] = 15'h7F37;
	tbl[1904] = 15'h7F39;
	tbl[1905] = 15'h7F3C;
	tbl[1906] = 15'h7F3F;
	tbl[1907] = 15'h7F42;
	tbl[1908] = 15'h7F44;
	tbl[1909] = 15'h7F47;
	tbl[1910] = 15'h7F4A;
	tbl[1911] = 15'h7F4C;
	tbl[1912] = 15'h7F4F;
	tbl[1913] = 15'h7F51;
	tbl[1914] = 15'h7F54;
	tbl[1915] = 15'h7F57;
	tbl[1916] = 15'h7F59;
	tbl[1917] = 15'h7F5C;
	tbl[1918] = 15'h7F5E;
	tbl[1919] = 15'h7F61;
	tbl[1920] = 15'h7F63;
	tbl[1921] = 15'h7F65;
	tbl[1922] = 15'h7F68;
	tbl[1923] = 15'h7F6A;
	tbl[1924] = 15'h7F6D;
	tbl[1925] = 15'h7F6F;
	tbl[1926] = 15'h7F71;
	tbl[1927] = 15'h7F74;
	tbl[1928] = 15'h7F76;
	tbl[1929] = 15'h7F78;
	tbl[1930] = 15'h7F7B;
	tbl[1931] = 15'h7F7D;
	tbl[1932] = 15'h7F7F;
	tbl[1933] = 15'h7F81;
	tbl[1934] = 15'h7F83;
	tbl[1935] = 15'h7F86;
	tbl[1936] = 15'h7F88;
	tbl[1937] = 15'h7F8A;
	tbl[1938] = 15'h7F8C;
	tbl[1939] = 15'h7F8E;
	tbl[1940] = 15'h7F90;
	tbl[1941] = 15'h7F92;
	tbl[1942] = 15'h7F94;
	tbl[1943] = 15'h7F96;
	tbl[1944] = 15'h7F98;
	tbl[1945] = 15'h7F9A;
	tbl[1946] = 15'h7F9C;
	tbl[1947] = 15'h7F9E;
	tbl[1948] = 15'h7FA0;
	tbl[1949] = 15'h7FA2;
	tbl[1950] = 15'h7FA4;
	tbl[1951] = 15'h7FA6;
	tbl[1952] = 15'h7FA7;
	tbl[1953] = 15'h7FA9;
	tbl[1954] = 15'h7FAB;
	tbl[1955] = 15'h7FAD;
	tbl[1956] = 15'h7FAF;
	tbl[1957] = 15'h7FB0;
	tbl[1958] = 15'h7FB2;
	tbl[1959] = 15'h7FB4;
	tbl[1960] = 15'h7FB6;
	tbl[1961] = 15'h7FB7;
	tbl[1962] = 15'h7FB9;
	tbl[1963] = 15'h7FBA;
	tbl[1964] = 15'h7FBC;
	tbl[1965] = 15'h7FBE;
	tbl[1966] = 15'h7FBF;
	tbl[1967] = 15'h7FC1;
	tbl[1968] = 15'h7FC2;
	tbl[1969] = 15'h7FC4;
	tbl[1970] = 15'h7FC5;
	tbl[1971] = 15'h7FC7;
	tbl[1972] = 15'h7FC8;
	tbl[1973] = 15'h7FCA;
	tbl[1974] = 15'h7FCB;
	tbl[1975] = 15'h7FCD;
	tbl[1976] = 15'h7FCE;
	tbl[1977] = 15'h7FCF;
	tbl[1978] = 15'h7FD1;
	tbl[1979] = 15'h7FD2;
	tbl[1980] = 15'h7FD3;
	tbl[1981] = 15'h7FD4;
	tbl[1982] = 15'h7FD6;
	tbl[1983] = 15'h7FD7;
	tbl[1984] = 15'h7FD8;
	tbl[1985] = 15'h7FD9;
	tbl[1986] = 15'h7FDB;
	tbl[1987] = 15'h7FDC;
	tbl[1988] = 15'h7FDD;
	tbl[1989] = 15'h7FDE;
	tbl[1990] = 15'h7FDF;
	tbl[1991] = 15'h7FE0;
	tbl[1992] = 15'h7FE1;
	tbl[1993] = 15'h7FE2;
	tbl[1994] = 15'h7FE3;
	tbl[1995] = 15'h7FE4;
	tbl[1996] = 15'h7FE5;
	tbl[1997] = 15'h7FE6;
	tbl[1998] = 15'h7FE7;
	tbl[1999] = 15'h7FE8;
	tbl[2000] = 15'h7FE9;
	tbl[2001] = 15'h7FEA;
	tbl[2002] = 15'h7FEB;
	tbl[2003] = 15'h7FEC;
	tbl[2004] = 15'h7FED;
	tbl[2005] = 15'h7FED;
	tbl[2006] = 15'h7FEE;
	tbl[2007] = 15'h7FEF;
	tbl[2008] = 15'h7FF0;
	tbl[2009] = 15'h7FF1;
	tbl[2010] = 15'h7FF1;
	tbl[2011] = 15'h7FF2;
	tbl[2012] = 15'h7FF3;
	tbl[2013] = 15'h7FF3;
	tbl[2014] = 15'h7FF4;
	tbl[2015] = 15'h7FF5;
	tbl[2016] = 15'h7FF5;
	tbl[2017] = 15'h7FF6;
	tbl[2018] = 15'h7FF6;
	tbl[2019] = 15'h7FF7;
	tbl[2020] = 15'h7FF7;
	tbl[2021] = 15'h7FF8;
	tbl[2022] = 15'h7FF8;
	tbl[2023] = 15'h7FF9;
	tbl[2024] = 15'h7FF9;
	tbl[2025] = 15'h7FFA;
	tbl[2026] = 15'h7FFA;
	tbl[2027] = 15'h7FFB;
	tbl[2028] = 15'h7FFB;
	tbl[2029] = 15'h7FFB;
	tbl[2030] = 15'h7FFC;
	tbl[2031] = 15'h7FFC;
	tbl[2032] = 15'h7FFC;
	tbl[2033] = 15'h7FFD;
	tbl[2034] = 15'h7FFD;
	tbl[2035] = 15'h7FFD;
	tbl[2036] = 15'h7FFD;
	tbl[2037] = 15'h7FFE;
	tbl[2038] = 15'h7FFE;
	tbl[2039] = 15'h7FFE;
	tbl[2040] = 15'h7FFE;
	tbl[2041] = 15'h7FFE;
	tbl[2042] = 15'h7FFE;
	tbl[2043] = 15'h7FFE;
	tbl[2044] = 15'h7FFE;
	tbl[2045] = 15'h7FFE;
	tbl[2046] = 15'h7FFE;
	tbl[2047] = 15'h7FFF;
end

endmodule
